	`define PADDR 32
	`define Reg_width 64
	`define USERSPACE 0
	`define Addr_space 17 
	`define byte_offset 2
	`define RV64 
